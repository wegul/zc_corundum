module moduleName (
    input  [2:0] iaa,
    output [0:0] baa
);

endmodule
